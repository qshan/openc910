/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @22
module ct_fadd_close_s1_d(
  close_adder0,
  close_adder1,
  close_op_chg,
  close_sum,
  ex1_double,
  ex1_single,
  ff1_pred,
  ff1_pred_onehot
);

// &Ports; @23
input   [53:0]  close_adder0;
input   [53:0]  close_adder1;
input           ex1_double;
input           ex1_single;
output          close_op_chg;
output  [53:0]  close_sum;
output  [5 :0]  ff1_pred;
output  [53:0]  ff1_pred_onehot;

// &Regs; @24
reg     [5 :0]  ff1_pred_t0;
reg     [53:0]  ff1_pred_t0_onehot;

// &Wires; @25
wire    [53:0]  close_adder0;
wire    [53:0]  close_adder0_t0;
wire    [53:0]  close_adder1;
wire    [53:0]  close_adder1_t0;
wire    [53:0]  close_ff1_a_t0;
wire    [53:0]  close_ff1_b_t0;
wire    [53:0]  close_ff1_c_t0;
wire    [53:0]  close_ff1_f_t0;
wire    [53:0]  close_ff1_g_t0;
wire    [53:0]  close_ff1_t_t0;
wire    [53:0]  close_ff1_z_t0;
wire    [53:0]  close_m1_oper2;
wire            close_op_chg;
wire    [53:0]  close_sum;
wire    [53:0]  close_sum_t0;
wire            ex1_double;
wire            ex1_single;
wire    [5 :0]  ff1_pred;
wire    [53:0]  ff1_pred_onehot;


//Three Type
//t0 : !src0_e_is_0 && !src1_e_is_0
//t1 : !src0_e_is_0 &&  src1_e_is_0
//t2 :  src0_e_is_0 &&  src1_e_is_0
//assign type0_sel = !src0_e_is_0 && !src1_e_is_0;
//assign type1_sel = !src0_e_is_0 &&  src1_e_is_0;
//assign type2_sel =  src0_e_is_0 &&  src1_e_is_0;

//assign close_sum[53:0]    = {54{type0_sel}} & close_sum_t0[53:0] |
//                            {54{type1_sel}} & close_sum_t1[53:0] |
//                            {54{type2_sel}} & close_sum_t2[53:0];
//assign close_sum_m1[53:0] = {54{type0_sel}} & close_sum_m1_t0[53:0] |
//                            {54{type1_sel}} & close_sum_m1_t1[53:0] |
//                            {54{type2_sel}} & close_sum_m1_t2[53:0];
//assign ff1_pred[53:0]     = {54{type0_sel}} & ff1_pred_t0_onehot[53:0] |
//                            {54{type1_sel}} & ff1_pred_t1_onehot[53:0] |
//                            {54{type2_sel}} & ff1_pred_t2[53:0];

assign close_sum[53:0]       = close_sum_t0[53:0];
//assign close_sum_m1[53:0]    = close_sum_m1_t0[53:0];
assign ff1_pred_onehot[53:0] = ff1_pred_t0_onehot[53:0];
assign ff1_pred[5:0]         = ff1_pred_t0[5:0];

assign close_op_chg       = close_sum[53];
// &Force("output","close_sum"); @51

assign close_adder0_t0[53:0] = close_adder0[53:0];
assign close_adder1_t0[53:0] = close_adder1[53:0];
//assign close_adder0_t1[53:0] = close_adder0[53:0];
//assign close_adder1_t1[53:0] = {1'b0, 1'b0, 22'b0, 29'b0};

assign close_m1_oper2[53:0]  = {54{ex1_double}} & 54'b10 |
                               {54{ex1_single}} & {24'b1,30'b0};
// &Force("nonport","close_sum_t0"); @60
// &Force("nonport","close_sum_m1_t0"); @61
// &Force("nonport","close_m1_oper2"); @62
//csky vperl_off
//close_sum0 for F0-F1
assign close_sum_t0[53:0] = $unsigned($signed(close_adder0_t0[53:0]) - $signed(close_adder1_t0[53:0]));
//close_sum0 for F1-F0
//close_sum select, keep sum not negative
//close_sum0_m1
//assign close_sum_m1_t0[53:0] = $unsigned($signed(close_adder0_t0[53:0])
//                                        - $signed(close_adder1_t0[53:0])
//                                        + $signed(close_m1_oper2[53:0]));
//csky vperl_on
//FF1 Logic of Close Path S0
//If predict first 1 set at r[n]
//Actual first 1 may set at r[n+1] or r[n]
//A and B are to oprand
assign close_ff1_a_t0[53:0] = close_adder0_t0[53:0];
assign close_ff1_b_t0[53:0] = close_adder1_t0[53:0];

//C = B && act_add || ~B && act_sub
assign close_ff1_c_t0[53:0] = ~close_ff1_b_t0[53:0];
//T = A^C  G=A&C  Z=(~A)&(~C)
assign close_ff1_t_t0[53:0] = close_ff1_a_t0[53:0] ^ close_ff1_c_t0[53:0];
assign close_ff1_g_t0[53:0] = close_ff1_a_t0[53:0] & close_ff1_c_t0[53:0];
assign close_ff1_z_t0[53:0] = (~close_ff1_a_t0[53:0]) & (~close_ff1_c_t0[53:0]);
//F :
//fn-1 = En[gi(~zi-1) + zi(~gi-1)] + (~En)[gi(~gi-1) + zi(~zi-1)], En=act_sub
//f0   = t1(g0En+z0) + (~t1)(z0En+g0)
//fi   = ti+1[gi(~zi-1) + zi(~gi-1)] + (~ti+1)[gi(~gi-1) + zi(~zi-1)]
assign close_ff1_f_t0[53]   =  ( close_ff1_g_t0[53] & (~close_ff1_z_t0[52])) |
                               ( close_ff1_z_t0[53] & (~close_ff1_g_t0[52]));
assign close_ff1_f_t0[0]    = (( close_ff1_t_t0[1]) & (close_ff1_g_t0[0] | close_ff1_z_t0[0])) |
                              ((~close_ff1_t_t0[1]) & (close_ff1_z_t0[0] | close_ff1_g_t0[0]));
assign close_ff1_f_t0[52:1] = (( close_ff1_t_t0[53:2]) & ((close_ff1_g_t0[52:1] & (~close_ff1_z_t0[51:0])) |
                               ( close_ff1_z_t0[52:1]  & (~close_ff1_g_t0[51:0]))))                     |
                              ((~close_ff1_t_t0[53:2]) & ((close_ff1_g_t0[52:1] & (~close_ff1_g_t0[51:0])) |
                               ( close_ff1_z_t0[52:1]  & (~close_ff1_z_t0[51:0]))));

// &CombBeg; @99
always @( close_ff1_f_t0[53:0])
begin
casez(close_ff1_f_t0[53:0])
  54'b1????_????????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b10000_00000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd0;
  end
  54'b01???_????????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b01000_00000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd1;
  end
  54'b001??_????????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00100_00000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd2;
  end
  54'b0001?_????????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00010_00000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd3;
  end
  54'b00001_????????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00001_00000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd4;
  end
  54'b00000_1???????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_10000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd5;
  end
  54'b00000_01??????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_01000000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd6;
  end
  54'b00000_001?????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00100000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd7;
  end
  54'b00000_0001????_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00010000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd8;
  end
  54'b00000_00001???_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00001000_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd9;
  end
  54'b00000_000001??_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000100_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd10;
  end
  54'b00000_0000001?_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000010_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd11;
  end
  54'b00000_00000001_????????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000001_00000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd12;
  end
  54'b00000_00000000_1???????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_10000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd13;
  end
  54'b00000_00000000_01??????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_01000000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd14;
  end
  54'b00000_00000000_001?????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00100000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd15;
  end
  54'b00000_00000000_0001????_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00010000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd16;
  end
  54'b00000_00000000_00001???_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00001000_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd17;
  end
  54'b00000_00000000_000001??_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000100_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd18;
  end
  54'b00000_00000000_0000001?_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000010_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd19;
  end
  54'b00000_00000000_00000001_????????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000001_00000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd20;
  end
  54'b00000_00000000_00000000_1???????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_10000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd21;
  end
  54'b00000_00000000_00000000_01??????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_01000000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd22;
  end
  54'b00000_00000000_00000000_001?????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00100000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd23;
  end
  54'b00000_00000000_00000000_0001????_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00010000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd24;
  end
  54'b00000_00000000_00000000_00001???_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00001000_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd25;
  end
  54'b00000_00000000_00000000_000001??_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000100_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd26;
  end
  54'b00000_00000000_00000000_0000001?_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000010_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd27;
  end
  54'b00000_00000000_00000000_00000001_????????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000001_00000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd28;
  end
  54'b00000_00000000_00000000_00000000_1???????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_10000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd29;
  end
  54'b00000_00000000_00000000_00000000_01??????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_01000000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd30;
  end
  54'b00000_00000000_00000000_00000000_001?????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00100000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd31;
  end
  54'b00000_00000000_00000000_00000000_0001????_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00010000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd32;
  end
  54'b00000_00000000_00000000_00000000_00001???_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00001000_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd33;
  end
  54'b00000_00000000_00000000_00000000_000001??_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000100_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd34;
  end
  54'b00000_00000000_00000000_00000000_0000001?_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000010_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd35;
  end
  54'b00000_00000000_00000000_00000000_00000001_????????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000001_00000000_000000000;
    ff1_pred_t0[5:0]         = 6'd36;
  end
  54'b00000_00000000_00000000_00000000_00000000_1???????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_10000000_000000000;
    ff1_pred_t0[5:0]         = 6'd37;
  end
  54'b00000_00000000_00000000_00000000_00000000_01??????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_01000000_000000000;
    ff1_pred_t0[5:0]         = 6'd38;
  end
  54'b00000_00000000_00000000_00000000_00000000_001?????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00100000_000000000;
    ff1_pred_t0[5:0]         = 6'd39;
  end
  54'b00000_00000000_00000000_00000000_00000000_0001????_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00010000_000000000;
    ff1_pred_t0[5:0]         = 6'd40;
  end
  54'b00000_00000000_00000000_00000000_00000000_00001???_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00001000_000000000;
    ff1_pred_t0[5:0]         = 6'd41;
  end
  54'b00000_00000000_00000000_00000000_00000000_000001??_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000100_000000000;
    ff1_pred_t0[5:0]         = 6'd42;
  end
  54'b00000_00000000_00000000_00000000_00000000_0000001?_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000010_000000000;
    ff1_pred_t0[5:0]         = 6'd43;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000001_????????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000001_000000000;
    ff1_pred_t0[5:0]         = 6'd44;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_1???????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_100000000;
    ff1_pred_t0[5:0]         = 6'd45;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_01??????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_010000000;
    ff1_pred_t0[5:0]         = 6'd46;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_001?????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_001000000;
    ff1_pred_t0[5:0]         = 6'd47;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_0001????? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000100000;
    ff1_pred_t0[5:0]         = 6'd48;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_00001???? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000010000;
    ff1_pred_t0[5:0]         = 6'd49;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_000001??? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000001000;
    ff1_pred_t0[5:0]         = 6'd50;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_0000001?? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000000100;
    ff1_pred_t0[5:0]         = 6'd51;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_00000001? : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000000010;
    ff1_pred_t0[5:0]         = 6'd52;
  end
  54'b00000_00000000_00000000_00000000_00000000_00000000_000000001 : begin
    ff1_pred_t0_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000000001;
    ff1_pred_t0[5:0]         = 6'd53;
  end

  default : begin
    ff1_pred_t0_onehot[53:0] = {54{1'bx}};
    ff1_pred_t0[5:0]         = {6{1'bx}};
  end
endcase
// &CombEnd; @323
end

////close_sum0 for F0-F1
//assign close_sum_t1[53:0] = close_adder0_t1[53:0] + ~close_adder1_t1[53:0] + 54'b1;
////close_sum0 for F1-F0
////close_sum select, keep sum not negative
////close_sum0_m1
//assign close_sum_m1_t1[53:0] = close_adder0_t1[53:0] + ~close_adder1_t1[53:0];
//
////FF1 Logic of Close Path S0
////If predict first 1 set at r[n]
////Actual first 1 may set at r[n+1] or r[n]
////A and B are to oprand
//assign close_ff1_a_t1[53:0] = close_adder0_t1[53:0];
//assign close_ff1_b_t1[53:0] = close_adder1_t1[53:0];
//
////C = B && act_add || ~B && act_sub
//assign close_ff1_c_t1[53:0] = ~close_ff1_b_t1[53:0];
////T = A^C  G=A&C  Z=(~A)&(~C)
//assign close_ff1_t_t1[53:0] = close_ff1_a_t1[53:0] ^ close_ff1_c_t1[53:0];
//assign close_ff1_g_t1[53:0] = close_ff1_a_t1[53:0] & close_ff1_c_t1[53:0];
//assign close_ff1_z_t1[53:0] = (~close_ff1_a_t1[53:0]) & (~close_ff1_c_t1[53:0]);
////F :
////fn-1 = En[gi(~zi-1) + zi(~gi-1)] + (~En)[gi(~gi-1) + zi(~zi-1)], En=act_sub
////f0   = t1(g0En+z0) + (~t1)(z0En+g0)
////fi   = ti+1[gi(~zi-1) + zi(~gi-1)] + (~ti+1)[gi(~gi-1) + zi(~zi-1)]
//assign close_ff1_f_t1[53]   =  ( close_ff1_g_t1[53] & (~close_ff1_z_t1[52])) |
//                               ( close_ff1_z_t1[53] & (~close_ff1_g_t1[52]));
//assign close_ff1_f_t1[0]    = (( close_ff1_t_t1[1]) & (close_ff1_g_t1[0] | close_ff1_z_t1[0])) |
//                              ((~close_ff1_t_t1[1]) & (close_ff1_z_t1[0] | close_ff1_g_t1[0]));
//assign close_ff1_f_t1[52:1] = (( close_ff1_t_t1[53:2]) & ((close_ff1_g_t1[52:1] & (~close_ff1_z_t1[51:0])) |
//                               ( close_ff1_z_t1[52:1]  & (~close_ff1_g_t1[51:0]))))                        |
//                              ((~close_ff1_t_t1[53:2]) & ((close_ff1_g_t1[52:1] & (~close_ff1_g_t1[51:0])) |
//                               ( close_ff1_z_t1[52:1]  & (~close_ff1_z_t1[51:0]))));
//
//
//&CombBeg;
//casez(close_ff1_f_t1[53:0])
//  54'b1????_????????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b10000_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd0;
//  end
//  54'b01???_????????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b01000_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd1;
//  end
//  54'b001??_????????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00100_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd2;
//  end
//  54'b0001?_????????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00010_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd3;
//  end
//  54'b00001_????????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00001_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd4;
//  end
//  54'b00000_1???????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_10000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd5;
//  end
//  54'b00000_01??????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_01000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd6;
//  end
//  54'b00000_001?????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00100000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd7;
//  end
//  54'b00000_0001????_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00010000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd8;
//  end
//  54'b00000_00001???_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00001000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd9;
//  end
//  54'b00000_000001??_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000100_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd10;
//  end
//  54'b00000_0000001?_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000010_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd11;
//  end
//  54'b00000_00000001_????????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000001_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd12;
//  end
//  54'b00000_00000000_1???????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_10000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd13;
//  end
//  54'b00000_00000000_01??????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_01000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd14;
//  end
//  54'b00000_00000000_001?????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00100000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd15;
//  end
//  54'b00000_00000000_0001????_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00010000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd16;
//  end
//  54'b00000_00000000_00001???_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00001000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd17;
//  end
//  54'b00000_00000000_000001??_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000100_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd18;
//  end
//  54'b00000_00000000_0000001?_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000010_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd19;
//  end
//  54'b00000_00000000_00000001_????????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000001_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd20;
//  end
//  54'b00000_00000000_00000000_1???????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_10000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd21;
//  end
//  54'b00000_00000000_00000000_01??????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_01000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd22;
//  end
//  54'b00000_00000000_00000000_001?????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00100000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd23;
//  end
//  54'b00000_00000000_00000000_0001????_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00010000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd24;
//  end
//  54'b00000_00000000_00000000_00001???_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00001000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd25;
//  end
//  54'b00000_00000000_00000000_000001??_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000100_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd26;
//  end
//  54'b00000_00000000_00000000_0000001?_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000010_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd27;
//  end
//  54'b00000_00000000_00000000_00000001_????????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000001_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd28;
//  end
//  54'b00000_00000000_00000000_00000000_1???????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_10000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd29;
//  end
//  54'b00000_00000000_00000000_00000000_01??????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_01000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd30;
//  end
//  54'b00000_00000000_00000000_00000000_001?????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00100000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd31;
//  end
//  54'b00000_00000000_00000000_00000000_0001????_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00010000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd32;
//  end
//  54'b00000_00000000_00000000_00000000_00001???_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00001000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd33;
//  end
//  54'b00000_00000000_00000000_00000000_000001??_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000100_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd34;
//  end
//  54'b00000_00000000_00000000_00000000_0000001?_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000010_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd35;
//  end
//  54'b00000_00000000_00000000_00000000_00000001_????????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000001_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd36;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_1???????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_10000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd37;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_01??????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_01000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd38;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_001?????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00100000_000000000;
//    ff1_pred_t1[5:0]         = 6'd39;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_0001????_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00010000_000000000;
//    ff1_pred_t1[5:0]         = 6'd40;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00001???_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00001000_000000000;
//    ff1_pred_t1[5:0]         = 6'd41;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_000001??_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000100_000000000;
//    ff1_pred_t1[5:0]         = 6'd42;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_0000001?_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000010_000000000;
//    ff1_pred_t1[5:0]         = 6'd43;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000001_????????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000001_000000000;
//    ff1_pred_t1[5:0]         = 6'd44;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_1???????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_100000000;
//    ff1_pred_t1[5:0]         = 6'd45;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_01??????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_010000000;
//    ff1_pred_t1[5:0]         = 6'd46;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_001?????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_001000000;
//    ff1_pred_t1[5:0]         = 6'd47;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_0001????? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000100000;
//    ff1_pred_t1[5:0]         = 6'd48;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_00001???? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000010000;
//    ff1_pred_t1[5:0]         = 6'd49;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_000001?? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000001000;
//    ff1_pred_t1[5:0]         = 6'd51;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_0000001? : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_00000010;
//    ff1_pred_t1[5:0]         = 6'd52;
//  end
//  54'b00000_00000000_00000000_00000000_00000000_00000000_00000001 : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_00000001;
//    ff1_pred_t1[5:0]         = 6'd53;
//  end
//  default : begin
//    ff1_pred_t1_onehot[53:0] = 54'b00000_00000000_00000000_00000000_00000000_00000000_000000000;
//    ff1_pred_t1[5:0]         = 6'd0;
//  end
//endcase
//&CombEnd;
//
//
//assign close_sum_t2[53:0]       = 54'b0;
//assign close_sum_m1_t2[53:0]    = 54'h1f_ffff_ffff_ffff;
//assign ff1_pred_t2_onehot[53:0] = 54'b0;
//assign ff1_pred_t2[5:0]         = 6'h0;
//
// &ModuleEnd; @586
endmodule



/*Copyright 2019-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

module compressor_32(a,b,c,s,ca);
parameter B_SIZE = 8;
input  [B_SIZE-1:0] a;
input  [B_SIZE-1:0] b;
input  [B_SIZE-1:0] c;
output [B_SIZE-1:0] s;
output [B_SIZE-1:0] ca;

wire [B_SIZE-1:0] s;
wire [B_SIZE-1:0]ca;

assign s[B_SIZE-1:0]  = a[B_SIZE-1:0]^b[B_SIZE-1:0]^c[B_SIZE-1:0];
assign ca[B_SIZE-1:0] = (a[B_SIZE-1:0]&b[B_SIZE-1:0])
                      | (c[B_SIZE-1:0]&b[B_SIZE-1:0])
                      | (a[B_SIZE-1:0]&c[B_SIZE-1:0]);

//reg   [B_SIZE-1:0]s,ca;
//integer i;
//always @(a[B_SIZE-1:0]
//      or b[B_SIZE-1:0]
//      or c[B_SIZE-1:0])
//begin
//  for(i= 0;i<B_SIZE;i=i+1) begin
//    {ca[i],s[i]} =  a[i] + b[i] +  c[i];
//  end
//end
endmodule
